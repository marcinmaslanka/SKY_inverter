magic
tech sky130A
timestamp 1737404755
<< nwell >>
rect 440 250 675 390
<< nmos >>
rect 580 115 595 215
<< pmos >>
rect 580 270 595 370
<< ndiff >>
rect 520 200 580 215
rect 520 130 535 200
rect 565 130 580 200
rect 520 115 580 130
rect 595 200 655 215
rect 595 130 610 200
rect 640 130 655 200
rect 595 115 655 130
<< pdiff >>
rect 520 355 580 370
rect 520 285 535 355
rect 565 285 580 355
rect 520 270 580 285
rect 595 355 655 370
rect 595 285 610 355
rect 640 285 655 355
rect 595 270 655 285
<< ndiffc >>
rect 535 130 565 200
rect 610 130 640 200
<< pdiffc >>
rect 535 285 565 355
rect 610 285 640 355
<< psubdiff >>
rect 460 200 520 215
rect 460 130 475 200
rect 505 130 520 200
rect 460 115 520 130
<< nsubdiff >>
rect 460 355 520 370
rect 460 285 475 355
rect 505 285 520 355
rect 460 270 520 285
<< psubdiffcont >>
rect 475 130 505 200
<< nsubdiffcont >>
rect 475 285 505 355
<< poly >>
rect 580 370 595 385
rect 580 215 595 270
rect 580 100 595 115
rect 555 90 595 100
rect 555 70 565 90
rect 585 70 595 90
rect 555 60 595 70
<< polycont >>
rect 565 70 585 90
<< locali >>
rect 465 355 575 365
rect 465 285 475 355
rect 505 285 535 355
rect 565 285 575 355
rect 465 275 575 285
rect 600 355 650 365
rect 600 285 610 355
rect 640 285 650 355
rect 600 275 650 285
rect 630 210 650 275
rect 465 200 575 210
rect 465 130 475 200
rect 505 130 535 200
rect 565 130 575 200
rect 465 120 575 130
rect 600 200 650 210
rect 600 130 610 200
rect 640 130 650 200
rect 600 120 650 130
rect 630 100 650 120
rect 440 90 595 100
rect 440 80 565 90
rect 555 70 565 80
rect 585 70 595 90
rect 630 80 675 100
rect 555 60 595 70
<< viali >>
rect 475 285 505 355
rect 535 285 565 355
rect 475 130 505 200
rect 535 130 565 200
<< metal1 >>
rect 440 355 675 365
rect 440 285 475 355
rect 505 285 535 355
rect 565 285 675 355
rect 440 275 675 285
rect 440 200 675 210
rect 440 130 475 200
rect 505 130 535 200
rect 565 130 675 200
rect 440 120 675 130
<< labels >>
rlabel locali 440 90 440 90 7 A
port 1 w
rlabel locali 675 90 675 90 3 Y
port 2 e
rlabel metal1 440 320 440 320 7 VP
port 3 w
rlabel metal1 440 165 440 165 7 VN
port 4 w
<< end >>
